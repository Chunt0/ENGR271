module parser (input logic [3:0] B, output logic [4:0] D);

    D[0] = B[0];
    D[1] = ;
    D[2] = ;
    D[3] = ;
    D[4] = ;
    
endmodule